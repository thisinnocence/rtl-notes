// xor_encryptor_tb.v (Corrected version 2)
`timescale 1ns / 1ps

module xor_encryptor_tb;

    // 信号声明和 DUT 实例化 (保持不变)
    reg  clk;
    reg  rst_n;
    reg  start;
    reg  [31:0] data_in;
    reg  [31:0] key_in;
    wire [31:0] data_out;
    wire done;

    xor_encryptor dut (
        .clk(clk),
        .rst_n(rst_n),
        .start(start),
        .data_in(data_in),
        .key_in(key_in),
        .data_out(data_out),
        .done(done)
    );

    initial begin
        clk = 1'b0;
        forever #5 clk = ~clk;
    end

    initial begin
        // 初始化
        rst_n = 1'b0;
        start = 1'b0;
        data_in = 32'hdeadbeef;
        key_in = 32'h12345678;

        // 1. 复位
        #10 rst_n = 1'b1;
        $display("----------------------------------------");
        $display("Test started.");

        // 2. 启动加密操作 (1个时钟周期)
        @(posedge clk);
        start = 1'b1;
        $display("Time=%0t, Starting encryption with:", $time);
        $display("Data_in  = 0x%h", data_in);
        $display("Key_in   = 0x%h", key_in);
        @(posedge clk);
        start = 1'b0;

        // 3. 等待状态机从 ENCRYPTING 到 DONE
        // 在这个时钟周期，done 信号会被置高
        @(posedge clk);
        
        // 4. 验证结果
        if (done) begin
            $display("Time=%0t, Encryption finished.", $time);
            $display("Expected output = 0x%h", data_in ^ key_in);
            $display("Actual output   = 0x%h", data_out);
            
            if (data_out == (data_in ^ key_in)) begin
                $display("----------------------------------------");
                $display("Test PASSED!");
                $display("----------------------------------------");
            end else begin
                $display("----------------------------------------");
                $display("Test FAILED: Incorrect output!");
                $display("----------------------------------------");
            end
        end else begin
            $display("Test FAILED: Done signal not received.");
        end

        // 5. 等待状态机从 DONE 回到 IDLE
        @(posedge clk);
        
        // 6. 再次运行
        data_in = 32'h01234567;
        key_in = 32'habcdef01;
        start = 1'b1;
        $display("----------------------------------------");
        $display("Test another case:");
        $display("Time=%0t, Starting encryption with:", $time);
        $display("Data_in  = 0x%h", data_in);
        $display("Key_in   = 0x%h", key_in);
        @(posedge clk);
        start = 1'b0;

        @(posedge clk);

        if (done && (data_out == (data_in ^ key_in))) begin
            $display("Time=%0t, Encryption finished.", $time);
            $display("Expected output = 0x%h", data_in ^ key_in);
            $display("Actual output   = 0x%h", data_out);
            $display("Test PASSED!");
        end else begin
            $display("Test FAILED!");
        end

        #10 $finish;
    end

endmodule